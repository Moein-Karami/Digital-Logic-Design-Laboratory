module TopDesign(input InFreq, ref_f, rst, adjust, start, input[3 :0]n, input [1 : 0]u, input [15 : 0]v,
		output done, output [20 : 0]exp_out);
	wire valid, acc_clk;

	FrequencyMultiplier fm(InFreq, ref_f, rst, adjust, n, acc_clk, valid);
	Wrapper wrapper(acc_clk, rst, start, , v, u, done, , , q, );
endmodule